`timescale 1ns / 1ps

module ALU(
	input clk,
	input rst,
	input [15:0] srcA,
	input [15:0] srcB,
	output [15:0] res,
	input [4:0] opsel,
	output ready,
	input [3:0] flags,
	output [3:0] flag_next
    );


endmodule
